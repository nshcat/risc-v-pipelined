module top(
    input logic clk_i,
    input logic rst_i
);

endmodule
