`ifndef _CORE_DEFINES_H
`define _CORE_DEFINES_H

// ======== Base data types ======== 
`define WORD_SIZE 32
typedef logic [`WORD_SIZE-1:0] word_t;

`endif